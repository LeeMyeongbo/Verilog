`timescale 1ns/1ps

module ALU_test(t1, t2, t3, p1);

output [7:0] t1, t2;
output [1:0] t3;
input  [7:0] p1;

reg [7:0] t1, t2;
reg [1:0] t3;

initial begin

    t1 <= 8'b0010_1011; t2 <= 8'b0001_1110;         // 덧셈 뺄셈 모두 정상 실행
    t3 <= 2'b00;
    #100;
    t3 <= 2'b01;
    #100;
    t3 <= 2'b10;
    #100;
    t3 <= 2'b11;

    #100;
    t1 <= 8'b1111_1001; t2 <= 8'b0101_1111;         // 덧셈 시 오버플로우 발생
    t3 <= 2'b00;
    #100;
    t3 <= 2'b01;
    #100;
    t3 <= 2'b10;
    #100;
    t3 <= 2'b11;

    #100;
    t1 <= 8'b0100_1011; t2 <= 8'b1000_0101;         // 뺄셈 시 오버플로우 발생
    t3 <= 2'b00;
    #100;
    t3 <= 2'b01;
    #100;
    t3 <= 2'b10;
    #100;
    t3 <= 2'b11;

    #100;
    $finish;
end

endmodule